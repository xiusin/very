module veb


pub interface AbstractBuilder<T>  {
}
