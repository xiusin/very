module dto

pub struct UserDto {
pub:
	username string [required]
	password string [required]
}
