module lark

pub struct AppAccessToken {
	code int
	msg string
	app_access_token string
	expire int
}