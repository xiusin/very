module contracts

pub interface Tabler {
	table_name() string
}
