module cache

fn test_di () ? {
	cache := new(Config{})?

	dump(cache)

}
