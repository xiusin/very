module builder

pub fn (builder &Builder) max(field string) ! {
}

pub fn (builder &Builder) min(field string) ! {
}

pub fn (builder &Builder) avg(field string) ! {
}

pub fn (builder &Builder) sum(field string) ! {
}

pub fn (builder &Builder) count(field string) ! {
}

pub fn (builder &Builder) value(field string) ! {
}

pub fn (builder &Builder) pluck(field string, index ...string) ! {
}
