module wechat

// 微信服务
enum WechatApiUrl {
	menu_create = '/cgi-bin/menu/create'
	menu_info = '/cgi-bin/get_current_selfmenu_info'
	menu_delete = '/cgi-bin/menu/delete'
	menu_get = '/cgi-bin/menu/get'
}
