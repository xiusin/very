module very

pub struct Request {
	http.Request
pub mut:
}
