module very

pub struct Request {
}
