module di

fn test_di() {
	println('hello')
}
