module builder

pub fn (b &Builder) max(field string) ! {
}

pub fn (b &Builder) min(field string) ! {
}

pub fn (b &Builder) avg(field string) ! {
}

pub fn (b &Builder) sum(field string) ! {
}

pub fn (b &Builder) count(field string) ! {
}

pub fn (b &Builder) value(field string) ! {
}

pub fn (b &Builder) pluck(field string, index ...string) ! {
}
