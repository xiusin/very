module builder

pub fn (builder &Builder) where_exists() {
}

pub fn (builder &Builder) or_where_exists() {
}

pub fn (builder &Builder) where_not_exists() {
}

pub fn (builder &Builder) or_where_not_exists() {
}
