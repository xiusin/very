module contracts
