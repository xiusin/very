module cache

struct Shard {
	hashmap map[u64]u32
}
