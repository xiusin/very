module di


pub struct Service {
	name string
mut:
 	instance voidptr
}
